/*
* @File name: Reservation_top
* @Author: Ruige Lee
* @Email: wut.ruigeli@gmail.com
* @Date:   2021-12-21 11:12:51
* @Last Modified by:   Ruige Lee
* @Last Modified time: 2021-12-21 11:39:13
*/


module Reservation_top(
  input         clock,
  input         reset
);


  wire   io_enq_0_ready;
  wire   io_enq_0_valid;
  wire  io_enq_0_bits_isa_fcsr_rw;


  wire    io_enq_1_ready;
  wire    io_enq_1_valid;
  wire    io_enq_1_bits_isa_fcsr_rs;
  wire    io_deq_0_ready;
  wire    io_deq_1_ready;

  wire       io_is_op_rsl_0_ready;
  wire       io_is_op_rsl_1_ready;
  wire       io_is_op_rsl_2_ready;
  wire       io_is_op_rsl_3_ready;

  wire io_is_wb_ack_0;
  wire io_is_wb_ack_1;
  wire io_is_wb_ack_2;


random_csr_req s_random_csr_req(
  .clock(clock),
  .reset(reset),

  .io_enq_0_ready(io_enq_0_ready),
  .io_enq_0_valid(io_enq_0_valid),
  .io_enq_0_bits_isa_fcsr_rw(io_enq_0_bits_isa_fcsr_rw),


  .io_enq_1_ready(io_enq_1_ready),
  .io_enq_1_valid(io_enq_1_valid),
  .io_enq_1_bits_isa_fcsr_rs(io_enq_1_bits_isa_fcsr_rs)


);

random_op_rsl s_random_op_rsl(
  .clock(clock),
  .reset(reset),

  .io_deq_0_ready(io_deq_0_ready),
  .io_deq_1_ready(io_deq_1_ready),

  .io_is_op_rsl_0_ready(io_is_op_rsl_0_ready),
  .io_is_op_rsl_1_ready(io_is_op_rsl_1_ready),
  .io_is_op_rsl_2_ready(io_is_op_rsl_2_ready),
  .io_is_op_rsl_3_ready(io_is_op_rsl_3_ready)

);


random_wb_ack s_random_wb_ack(

  .clock(clock),
  .reset(reset),

  .io_is_wb_ack_0(io_is_wb_ack_0),
  .io_is_wb_ack_1(io_is_wb_ack_1),
  .io_is_wb_ack_2(io_is_wb_ack_2)
);


Reservation_fpu s_Reservation_fpu(
  .clock(clock),
  .reset(reset),
  .io_enq_0_ready(io_enq_0_ready),
  .io_enq_0_valid(io_enq_0_valid),
  .io_enq_0_bits_isa_fmadd_s(1'b0),
  .io_enq_0_bits_isa_fmsub_s(1'b0),
  .io_enq_0_bits_isa_fnmsub_s(1'b0),
  .io_enq_0_bits_isa_fnmadd_s(1'b0),
  .io_enq_0_bits_isa_fadd_s(1'b0),
  .io_enq_0_bits_isa_fsub_s(1'b0),
  .io_enq_0_bits_isa_fmul_s(1'b0),
  .io_enq_0_bits_isa_fdiv_s(1'b0),
  .io_enq_0_bits_isa_fsqrt_s(1'b0),
  .io_enq_0_bits_isa_fsgnj_s(1'b0),
  .io_enq_0_bits_isa_fsgnjn_s(1'b0),
  .io_enq_0_bits_isa_fsgnjx_s(1'b0),
  .io_enq_0_bits_isa_fmin_s(1'b0),
  .io_enq_0_bits_isa_fmax_s(1'b0),
  .io_enq_0_bits_isa_fcvt_w_s(1'b0),
  .io_enq_0_bits_isa_fcvt_wu_s(1'b0),
  .io_enq_0_bits_isa_fmv_x_w(1'b0),
  .io_enq_0_bits_isa_feq_s(1'b0),
  .io_enq_0_bits_isa_flt_s(1'b0),
  .io_enq_0_bits_isa_fle_s(1'b0),
  .io_enq_0_bits_isa_fclass_s(1'b0),
  .io_enq_0_bits_isa_fcvt_s_w(1'b0),
  .io_enq_0_bits_isa_fcvt_s_wu(1'b0),
  .io_enq_0_bits_isa_fmv_w_x(1'b0),
  .io_enq_0_bits_isa_fcvt_l_s(1'b0),
  .io_enq_0_bits_isa_fcvt_lu_s(1'b0),
  .io_enq_0_bits_isa_fcvt_s_l(1'b0),
  .io_enq_0_bits_isa_fcvt_s_lu(1'b0),
  .io_enq_0_bits_isa_fmadd_d(1'b0),
  .io_enq_0_bits_isa_fmsub_d(1'b0),
  .io_enq_0_bits_isa_fnmsub_d(1'b0),
  .io_enq_0_bits_isa_fnmadd_d(1'b0),
  .io_enq_0_bits_isa_fadd_d(1'b0),
  .io_enq_0_bits_isa_fsub_d(1'b0),
  .io_enq_0_bits_isa_fmul_d(1'b0),
  .io_enq_0_bits_isa_fdiv_d(1'b0),
  .io_enq_0_bits_isa_fsqrt_d(1'b0),
  .io_enq_0_bits_isa_fsgnj_d(1'b0),
  .io_enq_0_bits_isa_fsgnjn_d(1'b0),
  .io_enq_0_bits_isa_fsgnjx_d(1'b0),
  .io_enq_0_bits_isa_fmin_d(1'b0),
  .io_enq_0_bits_isa_fmax_d(1'b0),
  .io_enq_0_bits_isa_fcvt_s_d(1'b0),
  .io_enq_0_bits_isa_fcvt_d_s(1'b0),
  .io_enq_0_bits_isa_feq_d(1'b0),
  .io_enq_0_bits_isa_flt_d(1'b0),
  .io_enq_0_bits_isa_fle_d(1'b0),
  .io_enq_0_bits_isa_fclass_d(1'b0),
  .io_enq_0_bits_isa_fcvt_w_d(1'b0),
  .io_enq_0_bits_isa_fcvt_wu_d(1'b0),
  .io_enq_0_bits_isa_fcvt_d_w(1'b0),
  .io_enq_0_bits_isa_fcvt_d_wu(1'b0),
  .io_enq_0_bits_isa_fcvt_l_d(1'b0),
  .io_enq_0_bits_isa_fcvt_lu_d(1'b0),
  .io_enq_0_bits_isa_fmv_x_d(1'b0),
  .io_enq_0_bits_isa_fcvt_d_l(1'b0),
  .io_enq_0_bits_isa_fcvt_d_lu(1'b0),
  .io_enq_0_bits_isa_fmv_d_x(1'b0),
  .io_enq_0_bits_isa_fcsr_rw(io_enq_0_bits_isa_fcsr_rw),
  .io_enq_0_bits_isa_fcsr_rs('d0),
  .io_enq_0_bits_isa_fcsr_rc('d0),
  .io_enq_0_bits_param_is_rvc('d0),
  .io_enq_0_bits_param_pc('d0),
  .io_enq_0_bits_param_imm('d0),
  .io_enq_0_bits_param_rm('d0),
  .io_enq_0_bits_param_rd0_raw('d0),
  .io_enq_0_bits_param_rs1_raw('d0),
  .io_enq_0_bits_param_rs2_raw('d0),
  .io_enq_0_bits_param_rs3_raw('d0),
  .io_enq_0_bits_phy_rd0('d0),
  .io_enq_0_bits_phy_rs1('d0),
  .io_enq_0_bits_phy_rs2('d0),
  .io_enq_0_bits_phy_rs3('d0),
  .io_enq_1_ready(io_enq_1_ready),
  .io_enq_1_valid(io_enq_1_valid),
  .io_enq_1_bits_isa_fmadd_s(1'b0),
  .io_enq_1_bits_isa_fmsub_s(1'b0),
  .io_enq_1_bits_isa_fnmsub_s(1'b0),
  .io_enq_1_bits_isa_fnmadd_s(1'b0),
  .io_enq_1_bits_isa_fadd_s(1'b0),
  .io_enq_1_bits_isa_fsub_s(1'b0),
  .io_enq_1_bits_isa_fmul_s(1'b0),
  .io_enq_1_bits_isa_fdiv_s(1'b0),
  .io_enq_1_bits_isa_fsqrt_s(1'b0),
  .io_enq_1_bits_isa_fsgnj_s(1'b0),
  .io_enq_1_bits_isa_fsgnjn_s(1'b0),
  .io_enq_1_bits_isa_fsgnjx_s(1'b0),
  .io_enq_1_bits_isa_fmin_s(1'b0),
  .io_enq_1_bits_isa_fmax_s(1'b0),
  .io_enq_1_bits_isa_fcvt_w_s(1'b0),
  .io_enq_1_bits_isa_fcvt_wu_s(1'b0),
  .io_enq_1_bits_isa_fmv_x_w(1'b0),
  .io_enq_1_bits_isa_feq_s(1'b0),
  .io_enq_1_bits_isa_flt_s(1'b0),
  .io_enq_1_bits_isa_fle_s(1'b0),
  .io_enq_1_bits_isa_fclass_s(1'b0),
  .io_enq_1_bits_isa_fcvt_s_w(1'b0),
  .io_enq_1_bits_isa_fcvt_s_wu(1'b0),
  .io_enq_1_bits_isa_fmv_w_x(1'b0),
  .io_enq_1_bits_isa_fcvt_l_s(1'b0),
  .io_enq_1_bits_isa_fcvt_lu_s(1'b0),
  .io_enq_1_bits_isa_fcvt_s_l(1'b0),
  .io_enq_1_bits_isa_fcvt_s_lu(1'b0),
  .io_enq_1_bits_isa_fmadd_d(1'b0),
  .io_enq_1_bits_isa_fmsub_d(1'b0),
  .io_enq_1_bits_isa_fnmsub_d(1'b0),
  .io_enq_1_bits_isa_fnmadd_d(1'b0),
  .io_enq_1_bits_isa_fadd_d(1'b0),
  .io_enq_1_bits_isa_fsub_d(1'b0),
  .io_enq_1_bits_isa_fmul_d(1'b0),
  .io_enq_1_bits_isa_fdiv_d(1'b0),
  .io_enq_1_bits_isa_fsqrt_d(1'b0),
  .io_enq_1_bits_isa_fsgnj_d(1'b0),
  .io_enq_1_bits_isa_fsgnjn_d(1'b0),
  .io_enq_1_bits_isa_fsgnjx_d(1'b0),
  .io_enq_1_bits_isa_fmin_d(1'b0),
  .io_enq_1_bits_isa_fmax_d(1'b0),
  .io_enq_1_bits_isa_fcvt_s_d(1'b0),
  .io_enq_1_bits_isa_fcvt_d_s(1'b0),
  .io_enq_1_bits_isa_feq_d(1'b0),
  .io_enq_1_bits_isa_flt_d(1'b0),
  .io_enq_1_bits_isa_fle_d(1'b0),
  .io_enq_1_bits_isa_fclass_d(1'b0),
  .io_enq_1_bits_isa_fcvt_w_d(1'b0),
  .io_enq_1_bits_isa_fcvt_wu_d(1'b0),
  .io_enq_1_bits_isa_fcvt_d_w(1'b0),
  .io_enq_1_bits_isa_fcvt_d_wu(1'b0),
  .io_enq_1_bits_isa_fcvt_l_d(1'b0),
  .io_enq_1_bits_isa_fcvt_lu_d(1'b0),
  .io_enq_1_bits_isa_fmv_x_d(1'b0),
  .io_enq_1_bits_isa_fcvt_d_l(1'b0),
  .io_enq_1_bits_isa_fcvt_d_lu(1'b0),
  .io_enq_1_bits_isa_fmv_d_x(1'b0),
  .io_enq_1_bits_isa_fcsr_rw(1'b0),
  .io_enq_1_bits_isa_fcsr_rs(io_enq_1_bits_isa_fcsr_rs),
  .io_enq_1_bits_isa_fcsr_rc('d0),
  .io_enq_1_bits_param_is_rvc('d0),
  .io_enq_1_bits_param_pc('d0),
  .io_enq_1_bits_param_imm('d0),
  .io_enq_1_bits_param_rm('d0),
  .io_enq_1_bits_param_rd0_raw('d0),
  .io_enq_1_bits_param_rs1_raw('d0),
  .io_enq_1_bits_param_rs2_raw('d0),
  .io_enq_1_bits_param_rs3_raw('d0),
  .io_enq_1_bits_phy_rd0('d0),
  .io_enq_1_bits_phy_rs1('d0),
  .io_enq_1_bits_phy_rs2('d0),
  .io_enq_1_bits_phy_rs3('d0),
  .io_deq_0_ready(io_deq_0_ready),
  .io_deq_0_valid(),
  .io_deq_0_bits_isa_fmadd_s(),
  .io_deq_0_bits_isa_fmsub_s(),
  .io_deq_0_bits_isa_fnmsub_s(),
  .io_deq_0_bits_isa_fnmadd_s(),
  .io_deq_0_bits_isa_fadd_s(),
  .io_deq_0_bits_isa_fsub_s(),
  .io_deq_0_bits_isa_fmul_s(),
  .io_deq_0_bits_isa_fdiv_s(),
  .io_deq_0_bits_isa_fsqrt_s(),
  .io_deq_0_bits_isa_fsgnj_s(),
  .io_deq_0_bits_isa_fsgnjn_s(),
  .io_deq_0_bits_isa_fsgnjx_s(),
  .io_deq_0_bits_isa_fmin_s(),
  .io_deq_0_bits_isa_fmax_s(),
  .io_deq_0_bits_isa_fcvt_w_s(),
  .io_deq_0_bits_isa_fcvt_wu_s(),
  .io_deq_0_bits_isa_fmv_x_w(),
  .io_deq_0_bits_isa_feq_s(),
  .io_deq_0_bits_isa_flt_s(),
  .io_deq_0_bits_isa_fle_s(),
  .io_deq_0_bits_isa_fclass_s(),
  .io_deq_0_bits_isa_fcvt_s_w(),
  .io_deq_0_bits_isa_fcvt_s_wu(),
  .io_deq_0_bits_isa_fmv_w_x(),
  .io_deq_0_bits_isa_fcvt_l_s(),
  .io_deq_0_bits_isa_fcvt_lu_s(),
  .io_deq_0_bits_isa_fcvt_s_l(),
  .io_deq_0_bits_isa_fcvt_s_lu(),
  .io_deq_0_bits_isa_fmadd_d(),
  .io_deq_0_bits_isa_fmsub_d(),
  .io_deq_0_bits_isa_fnmsub_d(),
  .io_deq_0_bits_isa_fnmadd_d(),
  .io_deq_0_bits_isa_fadd_d(),
  .io_deq_0_bits_isa_fsub_d(),
  .io_deq_0_bits_isa_fmul_d(),
  .io_deq_0_bits_isa_fdiv_d(),
  .io_deq_0_bits_isa_fsqrt_d(),
  .io_deq_0_bits_isa_fsgnj_d(),
  .io_deq_0_bits_isa_fsgnjn_d(),
  .io_deq_0_bits_isa_fsgnjx_d(),
  .io_deq_0_bits_isa_fmin_d(),
  .io_deq_0_bits_isa_fmax_d(),
  .io_deq_0_bits_isa_fcvt_s_d(),
  .io_deq_0_bits_isa_fcvt_d_s(),
  .io_deq_0_bits_isa_feq_d(),
  .io_deq_0_bits_isa_flt_d(),
  .io_deq_0_bits_isa_fle_d(),
  .io_deq_0_bits_isa_fclass_d(),
  .io_deq_0_bits_isa_fcvt_w_d(),
  .io_deq_0_bits_isa_fcvt_wu_d(),
  .io_deq_0_bits_isa_fcvt_d_w(),
  .io_deq_0_bits_isa_fcvt_d_wu(),
  .io_deq_0_bits_isa_fcvt_l_d(),
  .io_deq_0_bits_isa_fcvt_lu_d(),
  .io_deq_0_bits_isa_fmv_x_d(),
  .io_deq_0_bits_isa_fcvt_d_l(),
  .io_deq_0_bits_isa_fcvt_d_lu(),
  .io_deq_0_bits_isa_fmv_d_x(),
  .io_deq_0_bits_isa_fcsr_rw(),
  .io_deq_0_bits_isa_fcsr_rs(),
  .io_deq_0_bits_isa_fcsr_rc(),
  .io_deq_0_bits_param_is_rvc(),
  .io_deq_0_bits_param_pc(),
  .io_deq_0_bits_param_imm(),
  .io_deq_0_bits_param_rm(),
  .io_deq_0_bits_param_rd0_raw(),
  .io_deq_0_bits_param_rs1_raw(),
  .io_deq_0_bits_param_rs2_raw(),
  .io_deq_0_bits_param_rs3_raw(),
  .io_deq_0_bits_phy_rd0(),
  .io_deq_0_bits_phy_rs1(),
  .io_deq_0_bits_phy_rs2(),
  .io_deq_0_bits_phy_rs3(),
  .io_deq_1_ready(io_deq_1_ready),
  .io_deq_1_valid(),
  .io_deq_1_bits_isa_fmadd_s(),
  .io_deq_1_bits_isa_fmsub_s(),
  .io_deq_1_bits_isa_fnmsub_s(),
  .io_deq_1_bits_isa_fnmadd_s(),
  .io_deq_1_bits_isa_fadd_s(),
  .io_deq_1_bits_isa_fsub_s(),
  .io_deq_1_bits_isa_fmul_s(),
  .io_deq_1_bits_isa_fdiv_s(),
  .io_deq_1_bits_isa_fsqrt_s(),
  .io_deq_1_bits_isa_fsgnj_s(),
  .io_deq_1_bits_isa_fsgnjn_s(),
  .io_deq_1_bits_isa_fsgnjx_s(),
  .io_deq_1_bits_isa_fmin_s(),
  .io_deq_1_bits_isa_fmax_s(),
  .io_deq_1_bits_isa_fcvt_w_s(),
  .io_deq_1_bits_isa_fcvt_wu_s(),
  .io_deq_1_bits_isa_fmv_x_w(),
  .io_deq_1_bits_isa_feq_s(),
  .io_deq_1_bits_isa_flt_s(),
  .io_deq_1_bits_isa_fle_s(),
  .io_deq_1_bits_isa_fclass_s(),
  .io_deq_1_bits_isa_fcvt_s_w(),
  .io_deq_1_bits_isa_fcvt_s_wu(),
  .io_deq_1_bits_isa_fmv_w_x(),
  .io_deq_1_bits_isa_fcvt_l_s(),
  .io_deq_1_bits_isa_fcvt_lu_s(),
  .io_deq_1_bits_isa_fcvt_s_l(),
  .io_deq_1_bits_isa_fcvt_s_lu(),
  .io_deq_1_bits_isa_fmadd_d(),
  .io_deq_1_bits_isa_fmsub_d(),
  .io_deq_1_bits_isa_fnmsub_d(),
  .io_deq_1_bits_isa_fnmadd_d(),
  .io_deq_1_bits_isa_fadd_d(),
  .io_deq_1_bits_isa_fsub_d(),
  .io_deq_1_bits_isa_fmul_d(),
  .io_deq_1_bits_isa_fdiv_d(),
  .io_deq_1_bits_isa_fsqrt_d(),
  .io_deq_1_bits_isa_fsgnj_d(),
  .io_deq_1_bits_isa_fsgnjn_d(),
  .io_deq_1_bits_isa_fsgnjx_d(),
  .io_deq_1_bits_isa_fmin_d(),
  .io_deq_1_bits_isa_fmax_d(),
  .io_deq_1_bits_isa_fcvt_s_d(),
  .io_deq_1_bits_isa_fcvt_d_s(),
  .io_deq_1_bits_isa_feq_d(),
  .io_deq_1_bits_isa_flt_d(),
  .io_deq_1_bits_isa_fle_d(),
  .io_deq_1_bits_isa_fclass_d(),
  .io_deq_1_bits_isa_fcvt_w_d(),
  .io_deq_1_bits_isa_fcvt_wu_d(),
  .io_deq_1_bits_isa_fcvt_d_w(),
  .io_deq_1_bits_isa_fcvt_d_wu(),
  .io_deq_1_bits_isa_fcvt_l_d(),
  .io_deq_1_bits_isa_fcvt_lu_d(),
  .io_deq_1_bits_isa_fmv_x_d(),
  .io_deq_1_bits_isa_fcvt_d_l(),
  .io_deq_1_bits_isa_fcvt_d_lu(),
  .io_deq_1_bits_isa_fmv_d_x(),
  .io_deq_1_bits_isa_fcsr_rw(),
  .io_deq_1_bits_isa_fcsr_rs(),
  .io_deq_1_bits_isa_fcsr_rc(),
  .io_deq_1_bits_param_is_rvc(),
  .io_deq_1_bits_param_pc(),
  .io_deq_1_bits_param_imm(),
  .io_deq_1_bits_param_rm(),
  .io_deq_1_bits_param_rd0_raw(),
  .io_deq_1_bits_param_rs1_raw(),
  .io_deq_1_bits_param_rs2_raw(),
  .io_deq_1_bits_param_rs3_raw(),
  .io_deq_1_bits_phy_rd0(),
  .io_deq_1_bits_phy_rs1(),
  .io_deq_1_bits_phy_rs2(),
  .io_deq_1_bits_phy_rs3(),
  .io_is_op_rsl_0_ready(io_is_op_rsl_0_ready),
  .io_is_op_rsl_0_valid(),
  .io_is_op_rsl_0_bits_rd0(),
  .io_is_op_rsl_0_bits_rs1(),
  .io_is_op_rsl_0_bits_rs2(),
  .io_is_op_rsl_0_bits_rs3(),
  .io_is_op_rsl_1_ready(io_is_op_rsl_1_ready),
  .io_is_op_rsl_1_valid(),
  .io_is_op_rsl_1_bits_rd0(),
  .io_is_op_rsl_1_bits_rs1(),
  .io_is_op_rsl_1_bits_rs2(),
  .io_is_op_rsl_1_bits_rs3(),
  .io_is_op_rsl_2_ready(io_is_op_rsl_2_ready),
  .io_is_op_rsl_2_valid(),
  .io_is_op_rsl_2_bits_rd0(),
  .io_is_op_rsl_2_bits_rs1(),
  .io_is_op_rsl_2_bits_rs2(),
  .io_is_op_rsl_2_bits_rs3(),
  .io_is_op_rsl_3_ready(io_is_op_rsl_3_ready),
  .io_is_op_rsl_3_valid(),
  .io_is_op_rsl_3_bits_rd0(),
  .io_is_op_rsl_3_bits_rs1(),
  .io_is_op_rsl_3_bits_rs2(),
  .io_is_op_rsl_3_bits_rs3(),
  .io_is_wb_ack_0(io_is_wb_ack_0),
  .io_is_wb_ack_1(io_is_wb_ack_1),
  .io_is_wb_ack_2(io_is_wb_ack_2)
);



endmodule


